module seq_det_1011(
	input clk,rst,in,
	output reg out);

parameter S0=2'b00, S1=2'b01, S2=2'b10, S3=2'b11;

reg [1:0] cur_state, next_state;

always @(posedge clk or negedge rst)begin
	if(!rst)
		cur_state<= S0;
	else
		cur_state<= next_state;
end

always @(*) begin
	case(cur_state)
		S0: next_state= in? S1:S0;
		S1: next_state= in? S1:S2;
		S2: next_state= in? S3:S0;
		S3: next_state= in? S1:S2;
		default: next_state= S0;
	endcase
end

always @(*) begin
        out<=(cur_state==S3)&&(next_state==S1);
end

endmodule


